module InstructionMemory
#(parameter DATA_WIDTH=32, parameter ADDR_WIDTH=11)
(
	input [(DATA_WIDTH-1):0] data,
	input [(ADDR_WIDTH-1):0] read_addr, write_addr,
	input we, read_clock, write_clock,
	output reg [(DATA_WIDTH-1):0] q
);
	
	// Declare the RAM variable
	reg [DATA_WIDTH-1:0] ram[2**ADDR_WIDTH-1:0];
	
	initial 
	begin  
	ram[0] = 32'b01000100000000000000000000000000;//nop
ram[1] = 32'b01000100000000000000000000000000;//nop
ram[2] = 32'b00000100101011110000000000010100;//addi
ram[3] = 32'b00101100101011110000000000010011;//sw
ram[4] = 32'b00000100101011110000000000011000;//addi
ram[5] = 32'b00101100101011110000000000010111;//sw
ram[6] = 32'b00000100101011110000000000011100;//addi
ram[7] = 32'b00101100101011110000000000011011;//sw
ram[8] = 32'b00000100101011110000000000100000;//addi
ram[9] = 32'b00101100101011110000000000011111;//sw
ram[10] = 32'b00000100101011110000000000100100;//addi
ram[11] = 32'b00101100101011110000000000100011;//sw
ram[12] = 32'b10001100110000000000000010010111;//jump_reg
ram[13] = 32'b00101100011111110000000000000001;//sw
ram[14] = 32'b00000100010000100000000000000001;//addi
ram[15] = 32'b00000100010000100000000000000001;//addi
ram[16] = 32'b00101000101001110000000000011011;//lw
ram[17] = 32'b00101000011010000000000000000010;//lw
ram[18] = 32'b00000000111010000100100000000001;//add
ram[19] = 32'b00101001001001110000000000000000;//lw
ram[20] = 32'b00101100101001110000000000101011;//sw
ram[21] = 32'b00101000101001110000000000101011;//lw
ram[22] = 32'b00101000111001000000000000000000;//lw
ram[23] = 32'b00000100100100000000000000000000;//addi
ram[24] = 32'b00101000101001110000000000101011;//lw
ram[25] = 32'b00000100111010000000000000000010;//addi
ram[26] = 32'b00101001000001000000000000000000;//lw
ram[27] = 32'b00000100100100010000000000000000;//addi
ram[28] = 32'b00101000101001110000000000101011;//lw
ram[29] = 32'b00000100111010000000000000000011;//addi
ram[30] = 32'b00101001000001000000000000000000;//lw
ram[31] = 32'b00000100100100100000000000000000;//addi
ram[32] = 32'b00101000101001110000000000101011;//lw
ram[33] = 32'b00000100111010000000000000000100;//addi
ram[34] = 32'b00101001000001000000000000000000;//lw
ram[35] = 32'b00000100100100110000000000000000;//addi
ram[36] = 32'b00101000101001110000000000101011;//lw
ram[37] = 32'b00000100111010000000000000000101;//addi
ram[38] = 32'b00101001000001000000000000000000;//lw
ram[39] = 32'b00000100100101000000000000000000;//addi
ram[40] = 32'b00101000101001110000000000101011;//lw
ram[41] = 32'b00000100111010000000000000000110;//addi
ram[42] = 32'b00101001000001000000000000000000;//lw
ram[43] = 32'b00000100100101010000000000000000;//addi
ram[44] = 32'b00101000101001110000000000101011;//lw
ram[45] = 32'b00000100111010000000000000000111;//addi
ram[46] = 32'b00101001000001000000000000000000;//lw
ram[47] = 32'b00000100100101100000000000000000;//addi
ram[48] = 32'b00101000101001110000000000101011;//lw
ram[49] = 32'b00000100111010000000000000001000;//addi
ram[50] = 32'b00101001000001000000000000000000;//lw
ram[51] = 32'b00000100100101110000000000000000;//addi
ram[52] = 32'b00101000101001110000000000101011;//lw
ram[53] = 32'b00000100111010000000000000001001;//addi
ram[54] = 32'b00101001000001000000000000000000;//lw
ram[55] = 32'b00000100100110000000000000000000;//addi
ram[56] = 32'b00101000101001110000000000101011;//lw
ram[57] = 32'b00000100111010000000000000001010;//addi
ram[58] = 32'b00101001000001000000000000000000;//lw
ram[59] = 32'b00000100100110010000000000000000;//addi
ram[60] = 32'b00101000101001110000000000101011;//lw
ram[61] = 32'b00000100111010000000000000001011;//addi
ram[62] = 32'b00101001000001000000000000000000;//lw
ram[63] = 32'b00000100100110100000000000000000;//addi
ram[64] = 32'b00101000101001110000000000101011;//lw
ram[65] = 32'b00000100111010000000000000001100;//addi
ram[66] = 32'b00101001000001000000000000000000;//lw
ram[67] = 32'b00000100100110110000000000000000;//addi
ram[68] = 32'b00101000101001110000000000101011;//lw
ram[69] = 32'b00000100111010000000000000001101;//addi
ram[70] = 32'b00101001000001000000000000000000;//lw
ram[71] = 32'b00000100100111000000000000000000;//addi
ram[72] = 32'b00101000101001110000000000101011;//lw
ram[73] = 32'b00000100111010000000000000001110;//addi
ram[74] = 32'b00101001000001000000000000000000;//lw
ram[75] = 32'b00000100100111010000000000000000;//addi
ram[76] = 32'b00101000101001110000000000101011;//lw
ram[77] = 32'b00000100111010000000000000001111;//addi
ram[78] = 32'b00101001000001000000000000000000;//lw
ram[79] = 32'b00000100100111100000000000000000;//addi
ram[80] = 32'b00101000011111110000000000000001;//lw
ram[81] = 32'b00000011111000000000000000001100;//jr
ram[82] = 32'b00101100011111110000000000000001;//sw
ram[83] = 32'b00000100010000100000000000000001;//addi
ram[84] = 32'b00000100010000100000000000000001;//addi
ram[85] = 32'b00101000101001110000000000011011;//lw
ram[86] = 32'b00101000011010000000000000000010;//lw
ram[87] = 32'b00000000111010000100100000000001;//add
ram[88] = 32'b00101001001001110000000000000000;//lw
ram[89] = 32'b00101100101001110000000000101011;//sw
ram[90] = 32'b00000110000001000000000000000000;//addi
ram[91] = 32'b00101000101001110000000000101011;//lw
ram[92] = 32'b00101100111001000000000000000000;//sw
ram[93] = 32'b00000110001001000000000000000000;//addi
ram[94] = 32'b00101000101001110000000000101011;//lw
ram[95] = 32'b00000100111010000000000000000010;//addi
ram[96] = 32'b00101101000001000000000000000000;//sw
ram[97] = 32'b00000110010001000000000000000000;//addi
ram[98] = 32'b00101000101001110000000000101011;//lw
ram[99] = 32'b00000100111010000000000000000011;//addi
ram[100] = 32'b00101101000001000000000000000000;//sw
ram[101] = 32'b00000110011001000000000000000000;//addi
ram[102] = 32'b00101000101001110000000000101011;//lw
ram[103] = 32'b00000100111010000000000000000100;//addi
ram[104] = 32'b00101101000001000000000000000000;//sw
ram[105] = 32'b00000110100001000000000000000000;//addi
ram[106] = 32'b00101000101001110000000000101011;//lw
ram[107] = 32'b00000100111010000000000000000101;//addi
ram[108] = 32'b00101101000001000000000000000000;//sw
ram[109] = 32'b00000110101001000000000000000000;//addi
ram[110] = 32'b00101000101001110000000000101011;//lw
ram[111] = 32'b00000100111010000000000000000110;//addi
ram[112] = 32'b00101101000001000000000000000000;//sw
ram[113] = 32'b00000110110001000000000000000000;//addi
ram[114] = 32'b00101000101001110000000000101011;//lw
ram[115] = 32'b00000100111010000000000000000111;//addi
ram[116] = 32'b00101101000001000000000000000000;//sw
ram[117] = 32'b00000110111001000000000000000000;//addi
ram[118] = 32'b00101000101001110000000000101011;//lw
ram[119] = 32'b00000100111010000000000000001000;//addi
ram[120] = 32'b00101101000001000000000000000000;//sw
ram[121] = 32'b00000111000001000000000000000000;//addi
ram[122] = 32'b00101000101001110000000000101011;//lw
ram[123] = 32'b00000100111010000000000000001001;//addi
ram[124] = 32'b00101101000001000000000000000000;//sw
ram[125] = 32'b00000111001001000000000000000000;//addi
ram[126] = 32'b00101000101001110000000000101011;//lw
ram[127] = 32'b00000100111010000000000000001010;//addi
ram[128] = 32'b00101101000001000000000000000000;//sw
ram[129] = 32'b00000111010001000000000000000000;//addi
ram[130] = 32'b00101000101001110000000000101011;//lw
ram[131] = 32'b00000100111010000000000000001011;//addi
ram[132] = 32'b00101101000001000000000000000000;//sw
ram[133] = 32'b00000111011001000000000000000000;//addi
ram[134] = 32'b00101000101001110000000000101011;//lw
ram[135] = 32'b00000100111010000000000000001100;//addi
ram[136] = 32'b00101101000001000000000000000000;//sw
ram[137] = 32'b00000111100001000000000000000000;//addi
ram[138] = 32'b00101000101001110000000000101011;//lw
ram[139] = 32'b00000100111010000000000000001101;//addi
ram[140] = 32'b00101101000001000000000000000000;//sw
ram[141] = 32'b00000111101001000000000000000000;//addi
ram[142] = 32'b00101000101001110000000000101011;//lw
ram[143] = 32'b00000100111010000000000000001110;//addi
ram[144] = 32'b00101101000001000000000000000000;//sw
ram[145] = 32'b00000111110001000000000000000000;//addi
ram[146] = 32'b00101000101001110000000000101011;//lw
ram[147] = 32'b00000100111010000000000000001111;//addi
ram[148] = 32'b00101101000001000000000000000000;//sw
ram[149] = 32'b00101000011111110000000000000001;//lw
ram[150] = 32'b00000011111000000000000000001100;//jr
ram[151] = 32'b00000100000011110000000000000000;//addi
ram[152] = 32'b10010001111000000000000000000000;//show_pid
ram[153] = 32'b00101000101001110000000000010001;//lw
ram[154] = 32'b01100100111010000000000000000000;//seti
ram[155] = 32'b00011101000000000000000000010000;//beqz
ram[156] = 32'b00000100000011110000000000000000;//addi
ram[157] = 32'b00101100101011110000000000010000;//sw
ram[158] = 32'b00000100000011110000000000000001;//addi
ram[159] = 32'b00101100101011110000000000010001;//sw
ram[160] = 32'b00101000101001110000000000011111;//lw
ram[161] = 32'b00000100111010000000000000000000;//addi
ram[162] = 32'b00000100000011110000010000000000;//addi
ram[163] = 32'b00101101000011110000000000000000;//sw
ram[164] = 32'b00101000101001110000000000011111;//lw
ram[165] = 32'b00000100111010000000000000000001;//addi
ram[166] = 32'b00000100000011110000010100000000;//addi
ram[167] = 32'b00101101000011110000000000000000;//sw
ram[168] = 32'b00101000101001110000000000011111;//lw
ram[169] = 32'b00000100111010000000000000000010;//addi
ram[170] = 32'b00000100000011110000011000000000;//addi
ram[171] = 32'b00101101000011110000000000000000;//sw
ram[172] = 32'b00101000101001110000000000010000;//lw
ram[173] = 32'b01011000111010000000000000000000;//sgti
ram[174] = 32'b00011101000000000000000010000011;//beqz
ram[175] = 32'b00101000101001110000000000101100;//lw
ram[176] = 32'b01100100111010000000000000000001;//seti
ram[177] = 32'b00011101000000000000000000101100;//beqz
ram[178] = 32'b01101100100000000000000000000000;//get_pc
ram[179] = 32'b00101000101001110000000000010011;//lw
ram[180] = 32'b00101000101010000000000000010010;//lw
ram[181] = 32'b00000000111010000100100000000001;//add
ram[182] = 32'b00101101001001000000000000000000;//sw
ram[183] = 32'b00000111111001000000000000000000;//addi
ram[184] = 32'b00101100101001000000000000101110;//sw
ram[185] = 32'b00000110000001000000000000000000;//addi
ram[186] = 32'b00101000101001110000000000100011;//lw
ram[187] = 32'b00101000101010000000000000010010;//lw
ram[188] = 32'b00000000111010000100100000000001;//add
ram[189] = 32'b00101101001001000000000000000000;//sw
ram[190] = 32'b00101000101001110000000000100011;//lw
ram[191] = 32'b00101000101010000000000000010010;//lw
ram[192] = 32'b00000000111010000100100000000001;//add
ram[193] = 32'b00101001001001110000000000000000;//lw
ram[194] = 32'b01100100111010000000000000000000;//seti
ram[195] = 32'b00011101000000000000000000000100;//beqz
ram[196] = 32'b00101000101001110000000000010000;//lw
ram[197] = 32'b00000100111010001111111111111111;//addi
ram[198] = 32'b00101100101010000000000000010000;//sw
ram[199] = 32'b10001100110000000000000011011101;//jump_reg
ram[200] = 32'b00101000101001110000000000011011;//lw
ram[201] = 32'b00101000101010000000000000010010;//lw
ram[202] = 32'b00000000111010000100100000000001;//add
ram[203] = 32'b00101001001001110000000000000000;//lw
ram[204] = 32'b00000100111010000000000000000001;//addi
ram[205] = 32'b00101100101010000000000000101011;//sw
ram[206] = 32'b00101000101001110000000000101110;//lw
ram[207] = 32'b00101000101010000000000000101011;//lw
ram[208] = 32'b00101101000001110000000000000000;//sw
ram[209] = 32'b00101000101001110000000000010010;//lw
ram[210] = 32'b00101100010001110000000000000000;//sw
ram[211] = 32'b00000100010000100000000000000001;//addi
ram[212] = 32'b00101100010000110000000000000000;//sw
ram[213] = 32'b00000100010000110000000000000000;//addi
ram[214] = 32'b00000100010000100000000000000001;//addi
ram[215] = 32'b00101100011001110000000000000010;//sw
ram[216] = 32'b10001000110000000000000001010010;//jal_reg
ram[217] = 32'b00000100011000100000000000000000;//addi
ram[218] = 32'b00101000011000110000000000000000;//lw
ram[219] = 32'b00000100010000101111111111111111;//addi
ram[220] = 32'b00101000010001110000000000000000;//lw
ram[221] = 32'b10001100110000000000000011100110;//jump_reg
ram[222] = 32'b00101000101001110000000000100011;//lw
ram[223] = 32'b00101000101010000000000000010010;//lw
ram[224] = 32'b00000000111010000100100000000001;//add
ram[225] = 32'b00000100000011110000000000000000;//addi
ram[226] = 32'b00101101001011110000000000000000;//sw
ram[227] = 32'b00101000101001110000000000010000;//lw
ram[228] = 32'b00000100111010001111111111111111;//addi
ram[229] = 32'b00101100101010000000000000010000;//sw
ram[230] = 32'b00101000101001110000000000010000;//lw
ram[231] = 32'b01011000111010000000000000000000;//sgti
ram[232] = 32'b00011101000000000000000001000110;//beqz
ram[233] = 32'b00101000101001110000000000010010;//lw
ram[234] = 32'b00000100111010000000000000000001;//addi
ram[235] = 32'b00101100101010000000000000010010;//sw
ram[236] = 32'b00101000101001110000000000010010;//lw
ram[237] = 32'b01100100111010000000000000000011;//seti
ram[238] = 32'b00011101000000000000000000000010;//beqz
ram[239] = 32'b00000100000011110000000000000000;//addi
ram[240] = 32'b00101100101011110000000000010010;//sw
ram[241] = 32'b00101000101001110000000000100011;//lw
ram[242] = 32'b00101000101010000000000000010010;//lw
ram[243] = 32'b00000000111010000100100000000001;//add
ram[244] = 32'b00101001001001110000000000000000;//lw
ram[245] = 32'b01101000111010000000000000000001;//sdti
ram[246] = 32'b00011101000000000000000000001001;//beqz
ram[247] = 32'b00101000101001110000000000010010;//lw
ram[248] = 32'b00000100111010000000000000000001;//addi
ram[249] = 32'b00101100101010000000000000010010;//sw
ram[250] = 32'b00101000101001110000000000010010;//lw
ram[251] = 32'b01100100111010000000000000000011;//seti
ram[252] = 32'b00011101000000000000000000000010;//beqz
ram[253] = 32'b00000100000011110000000000000000;//addi
ram[254] = 32'b00101100101011110000000000010010;//sw
ram[255] = 32'b10001100110000000000000011110001;//jump_reg
ram[256] = 32'b00101000101001110000000000010010;//lw
ram[257] = 32'b00101100010001110000000000000000;//sw
ram[258] = 32'b00000100010000100000000000000001;//addi
ram[259] = 32'b00101100010000110000000000000000;//sw
ram[260] = 32'b00000100010000110000000000000000;//addi
ram[261] = 32'b00000100010000100000000000000001;//addi
ram[262] = 32'b00101100011001110000000000000010;//sw
ram[263] = 32'b10001000110000000000000000001101;//jal_reg
ram[264] = 32'b00000100011000100000000000000000;//addi
ram[265] = 32'b00101000011000110000000000000000;//lw
ram[266] = 32'b00000100010000101111111111111111;//addi
ram[267] = 32'b00101000010001110000000000000000;//lw
ram[268] = 32'b00101000101001110000000000011011;//lw
ram[269] = 32'b00101000101010000000000000010010;//lw
ram[270] = 32'b00000000111010000100100000000001;//add
ram[271] = 32'b00101001001001110000000000000000;//lw
ram[272] = 32'b00000100111010000000000000000001;//addi
ram[273] = 32'b00101100101010000000000000101011;//sw
ram[274] = 32'b00101000101001110000000000101011;//lw
ram[275] = 32'b00101000111001000000000000000000;//lw
ram[276] = 32'b00101100101001000000000000101010;//sw
ram[277] = 32'b00101000101001110000000000101010;//lw
ram[278] = 32'b00000100111111110000000000000000;//addi
ram[279] = 32'b00101000101001110000000000010000;//lw
ram[280] = 32'b01100100111010000000000000000001;//seti
ram[281] = 32'b00011101000000000000000000000010;//beqz
ram[282] = 32'b00000100000011110000000000000000;//addi
ram[283] = 32'b00101100101011110000000000101100;//sw
ram[284] = 32'b00101000101001110000000000010010;//lw
ram[285] = 32'b00000100111010000000000000000001;//addi
ram[286] = 32'b10010001000000000000000000000000;//show_pid
ram[287] = 32'b00101000101001110000000000101100;//lw
ram[288] = 32'b01100100111010000000000000000001;//seti
ram[289] = 32'b00011101000000000000000000000111;//beqz
ram[290] = 32'b00101000101001110000000000010011;//lw
ram[291] = 32'b00101000101010000000000000010010;//lw
ram[292] = 32'b00000000111010000100100000000001;//add
ram[293] = 32'b00101001001001110000000000000000;//lw
ram[294] = 32'b01110000000000000000000000000000;//enable_timer
ram[295] = 32'b00000000111000000000000000001100;//jr
ram[296] = 32'b10001100110000000000000100101110;//jump_reg
ram[297] = 32'b00101000101001110000000000010011;//lw
ram[298] = 32'b00101000101010000000000000010010;//lw
ram[299] = 32'b00000000111010000100100000000001;//add
ram[300] = 32'b00101001001001110000000000000000;//lw
ram[301] = 32'b00000000111000000000000000001100;//jr
ram[302] = 32'b10001100110000000000000100110001;//jump_reg
ram[303] = 32'b00000100000011110000001111100111;//addi
ram[304] = 32'b01010001111000000000000000000000;//output
ram[305] = 32'b10001100110000000000000111000010;//jump_reg
ram[306] = 32'b00000100000011110000000000000010;//addi
ram[307] = 32'b00101100101011110000000000010000;//sw
ram[308] = 32'b00000100000011110000000000000000;//addi
ram[309] = 32'b00101100101011110000000000101100;//sw
ram[310] = 32'b00000100000011110000000000000000;//addi
ram[311] = 32'b00101100101011110000000000101000;//sw
ram[312] = 32'b00101000101001110000000000101000;//lw
ram[313] = 32'b00101000101010000000000000010000;//lw
ram[314] = 32'b00000000111010000100100000001000;//slt
ram[315] = 32'b00011101001000000000000001011110;//beqz
ram[316] = 32'b00101000101001110000000000011111;//lw
ram[317] = 32'b00101000101010000000000000101000;//lw
ram[318] = 32'b00000000111010000100100000000001;//add
ram[319] = 32'b00101001001001110000000000000000;//lw
ram[320] = 32'b00101000101010000000000000010111;//lw
ram[321] = 32'b00101000101010010000000000101000;//lw
ram[322] = 32'b00000001000010010101000000000001;//add
ram[323] = 32'b00101101010001110000000000000000;//sw
ram[324] = 32'b00101000101001110000000000101000;//lw
ram[325] = 32'b00000100111010000000000000000001;//addi
ram[326] = 32'b00001001000001110000001000000000;//multi
ram[327] = 32'b00101000101010000000000000011011;//lw
ram[328] = 32'b00101000101010010000000000101000;//lw
ram[329] = 32'b00000001000010010101000000000001;//add
ram[330] = 32'b00101101010001110000000000000000;//sw
ram[331] = 32'b00101000101001110000000000011111;//lw
ram[332] = 32'b00101000101010000000000000101000;//lw
ram[333] = 32'b00000000111010000100100000000001;//add
ram[334] = 32'b00101001001001110000000000000000;//lw
ram[335] = 32'b00101000101010000000000000010011;//lw
ram[336] = 32'b00101000101010010000000000101000;//lw
ram[337] = 32'b00000001000010010101000000000001;//add
ram[338] = 32'b00101101010001110000000000000000;//sw
ram[339] = 32'b00101000101001110000000000100011;//lw
ram[340] = 32'b00101000101010000000000000101000;//lw
ram[341] = 32'b00000000111010000100100000000001;//add
ram[342] = 32'b00000100000011110000000000000001;//addi
ram[343] = 32'b00101101001011110000000000000000;//sw
ram[344] = 32'b00101000101001110000000000011011;//lw
ram[345] = 32'b00101000101010000000000000101000;//lw
ram[346] = 32'b00000000111010000100100000000001;//add
ram[347] = 32'b00101001001001110000000000000000;//lw
ram[348] = 32'b00000100111010000000000001000010;//addi
ram[349] = 32'b00101100101010000000000000101010;//sw
ram[350] = 32'b00101000101001110000000000011011;//lw
ram[351] = 32'b00101000101010000000000000101000;//lw
ram[352] = 32'b00000000111010000100100000000001;//add
ram[353] = 32'b00101001001001110000000000000000;//lw
ram[354] = 32'b00000100111010000000000000000010;//addi
ram[355] = 32'b00101100101010000000000000101011;//sw
ram[356] = 32'b00101000101001110000000000101010;//lw
ram[357] = 32'b00101000101010000000000000101011;//lw
ram[358] = 32'b00101101000001110000000000000000;//sw
ram[359] = 32'b00101000101001110000000000011011;//lw
ram[360] = 32'b00101000101010000000000000101000;//lw
ram[361] = 32'b00000000111010000100100000000001;//add
ram[362] = 32'b00101001001001110000000000000000;//lw
ram[363] = 32'b00000100111010000000000000000011;//addi
ram[364] = 32'b00101100101010000000000000101011;//sw
ram[365] = 32'b00101000101001110000000000101010;//lw
ram[366] = 32'b00101000101010000000000000101011;//lw
ram[367] = 32'b00101101000001110000000000000000;//sw
ram[368] = 32'b00101000101001110000000000011011;//lw
ram[369] = 32'b00101000101010000000000000101000;//lw
ram[370] = 32'b00000000111010000100100000000001;//add
ram[371] = 32'b00101001001001110000000000000000;//lw
ram[372] = 32'b00000100111010000000000000000101;//addi
ram[373] = 32'b00101100101010000000000000101011;//sw
ram[374] = 32'b00101000101001110000000000011011;//lw
ram[375] = 32'b00101000101010000000000000101000;//lw
ram[376] = 32'b00000000111010000100100000000001;//add
ram[377] = 32'b00101001001001110000000000000000;//lw
ram[378] = 32'b00101100101001110000000000101010;//sw
ram[379] = 32'b00101000101001110000000000101010;//lw
ram[380] = 32'b00101000101010000000000000101011;//lw
ram[381] = 32'b00101101000001110000000000000000;//sw
ram[382] = 32'b00101000101001110000000000011011;//lw
ram[383] = 32'b00101000101010000000000000101000;//lw
ram[384] = 32'b00000000111010000100100000000001;//add
ram[385] = 32'b00101001001001110000000000000000;//lw
ram[386] = 32'b00101100101001110000000000101011;//sw
ram[387] = 32'b00000100000011110000000000000001;//addi
ram[388] = 32'b00101100101011110000000000101010;//sw
ram[389] = 32'b00101000101001110000000000101010;//lw
ram[390] = 32'b00101000101010000000000000101011;//lw
ram[391] = 32'b00101101000001110000000000000000;//sw
ram[392] = 32'b00101000101001110000000000011011;//lw
ram[393] = 32'b00101000101010000000000000101000;//lw
ram[394] = 32'b00000000111010000100100000000001;//add
ram[395] = 32'b00101001001001110000000000000000;//lw
ram[396] = 32'b00000100111010000000000000000110;//addi
ram[397] = 32'b00101100101010000000000000101011;//sw
ram[398] = 32'b00101000101001110000000000010111;//lw
ram[399] = 32'b00101000101010000000000000101000;//lw
ram[400] = 32'b00000000111010000100100000000001;//add
ram[401] = 32'b00101001001001110000000000000000;//lw
ram[402] = 32'b00101100101001110000000000101010;//sw
ram[403] = 32'b00101000101001110000000000101010;//lw
ram[404] = 32'b00101000101010000000000000101011;//lw
ram[405] = 32'b00101101000001110000000000000000;//sw
ram[406] = 32'b00101000101001110000000000101000;//lw
ram[407] = 32'b00000100111010000000000000000001;//addi
ram[408] = 32'b00101100101010000000000000101000;//sw
ram[409] = 32'b10001100110000000000000100111000;//jump_reg
ram[410] = 32'b00000100000011110000000000000000;//addi
ram[411] = 32'b00101100101011110000000000010010;//sw
ram[412] = 32'b00101100010000110000000000000000;//sw
ram[413] = 32'b00000100010000110000000000000000;//addi
ram[414] = 32'b00000100010000100000000000000001;//addi
ram[415] = 32'b00000100000011110000000000000000;//addi
ram[416] = 32'b00101100011011110000000000000010;//sw
ram[417] = 32'b10001000110000000000000000001101;//jal_reg
ram[418] = 32'b00000100011000100000000000000000;//addi
ram[419] = 32'b00101000011000110000000000000000;//lw
ram[420] = 32'b00101000101001110000000000011011;//lw
ram[421] = 32'b00000100111010000000000000000000;//addi
ram[422] = 32'b00101001000001110000000000000000;//lw
ram[423] = 32'b00000100111010000000000000000001;//addi
ram[424] = 32'b00101100101010000000000000101011;//sw
ram[425] = 32'b00101000101001110000000000101011;//lw
ram[426] = 32'b00101000111001000000000000000000;//lw
ram[427] = 32'b00101100101001000000000000101010;//sw
ram[428] = 32'b00101000101001110000000000101010;//lw
ram[429] = 32'b00000100111111110000000000000000;//addi
ram[430] = 32'b00101000101001110000000000010000;//lw
ram[431] = 32'b01100100111010000000000000000001;//seti
ram[432] = 32'b00011101000000000000000000000010;//beqz
ram[433] = 32'b00000100000011110000000000000000;//addi
ram[434] = 32'b00101100101011110000000000101100;//sw
ram[435] = 32'b00000100000011110000000000000001;//addi
ram[436] = 32'b10010001111000000000000000000000;//show_pid
ram[437] = 32'b00101000101001110000000000101100;//lw
ram[438] = 32'b01100100111010000000000000000001;//seti
ram[439] = 32'b00011101000000000000000000000110;//beqz
ram[440] = 32'b00101000101001110000000000010011;//lw
ram[441] = 32'b00000100111010000000000000000000;//addi
ram[442] = 32'b00101001000001110000000000000000;//lw
ram[443] = 32'b01110000000000000000000000000000;//enable_timer
ram[444] = 32'b00000000111000000000000000001100;//jr
ram[445] = 32'b10001100110000000000000111000010;//jump_reg
ram[446] = 32'b00101000101001110000000000010011;//lw
ram[447] = 32'b00000100111010000000000000000000;//addi
ram[448] = 32'b00101001000001110000000000000000;//lw
ram[449] = 32'b00000000111000000000000000001100;//jr

	
	
//		ram[0] = 32'b01000100000000000000000000000000;//nop
//		ram[1] = 32'b01000100000000000000000000000000;//nop
//		ram[2] = 32'b00000100101011110000000000010100;//addi
//		ram[3] = 32'b00101100101011110000000000010011;//sw
//		ram[4] = 32'b00000100101011110000000000011000;//addi
//		ram[5] = 32'b00101100101011110000000000010111;//sw
//		ram[6] = 32'b00000100101011110000000000011100;//addi
//		ram[7] = 32'b00101100101011110000000000011011;//sw
//		ram[8] = 32'b00000100101011110000000000100000;//addi
//		ram[9] = 32'b00101100101011110000000000011111;//sw
//		ram[10] = 32'b00000100101011110000000000100100;//addi
//		ram[11] = 32'b00101100101011110000000000100011;//sw
//		ram[12] = 32'b10001100110000000000000010010111;//jump_reg
//		ram[13] = 32'b00101100011111110000000000000001;//sw
//		ram[14] = 32'b00000100010000100000000000000001;//addi
//		ram[15] = 32'b00000100010000100000000000000001;//addi
//		ram[16] = 32'b00101000101001110000000000011011;//lw
//		ram[17] = 32'b00101000011010000000000000000010;//lw
//		ram[18] = 32'b00000000111010000100100000000001;//add
//		ram[19] = 32'b00101001001001110000000000000000;//lw
//		ram[20] = 32'b00101100101001110000000000101011;//sw
//		ram[21] = 32'b00101000101001110000000000101011;//lw
//		ram[22] = 32'b00101000111001000000000000000000;//lw
//		ram[23] = 32'b00000100100100000000000000000000;//addi
//		ram[24] = 32'b00101000101001110000000000101011;//lw
//		ram[25] = 32'b00000100111010000000000000000010;//addi
//		ram[26] = 32'b00101001000001000000000000000000;//lw
//		ram[27] = 32'b00000100100100010000000000000000;//addi
//		ram[28] = 32'b00101000101001110000000000101011;//lw
//		ram[29] = 32'b00000100111010000000000000000011;//addi
//		ram[30] = 32'b00101001000001000000000000000000;//lw
//		ram[31] = 32'b00000100100100100000000000000000;//addi
//		ram[32] = 32'b00101000101001110000000000101011;//lw
//		ram[33] = 32'b00000100111010000000000000000100;//addi
//		ram[34] = 32'b00101001000001000000000000000000;//lw
//		ram[35] = 32'b00000100100100110000000000000000;//addi
//		ram[36] = 32'b00101000101001110000000000101011;//lw
//		ram[37] = 32'b00000100111010000000000000000101;//addi
//		ram[38] = 32'b00101001000001000000000000000000;//lw
//		ram[39] = 32'b00000100100101000000000000000000;//addi
//		ram[40] = 32'b00101000101001110000000000101011;//lw
//		ram[41] = 32'b00000100111010000000000000000110;//addi
//		ram[42] = 32'b00101001000001000000000000000000;//lw
//		ram[43] = 32'b00000100100101010000000000000000;//addi
//		ram[44] = 32'b00101000101001110000000000101011;//lw
//		ram[45] = 32'b00000100111010000000000000000111;//addi
//		ram[46] = 32'b00101001000001000000000000000000;//lw
//		ram[47] = 32'b00000100100101100000000000000000;//addi
//		ram[48] = 32'b00101000101001110000000000101011;//lw
//		ram[49] = 32'b00000100111010000000000000001000;//addi
//		ram[50] = 32'b00101001000001000000000000000000;//lw
//		ram[51] = 32'b00000100100101110000000000000000;//addi
//		ram[52] = 32'b00101000101001110000000000101011;//lw
//		ram[53] = 32'b00000100111010000000000000001001;//addi
//		ram[54] = 32'b00101001000001000000000000000000;//lw
//		ram[55] = 32'b00000100100110000000000000000000;//addi
//		ram[56] = 32'b00101000101001110000000000101011;//lw
//		ram[57] = 32'b00000100111010000000000000001010;//addi
//		ram[58] = 32'b00101001000001000000000000000000;//lw
//		ram[59] = 32'b00000100100110010000000000000000;//addi
//		ram[60] = 32'b00101000101001110000000000101011;//lw
//		ram[61] = 32'b00000100111010000000000000001011;//addi
//		ram[62] = 32'b00101001000001000000000000000000;//lw
//		ram[63] = 32'b00000100100110100000000000000000;//addi
//		ram[64] = 32'b00101000101001110000000000101011;//lw
//		ram[65] = 32'b00000100111010000000000000001100;//addi
//		ram[66] = 32'b00101001000001000000000000000000;//lw
//		ram[67] = 32'b00000100100110110000000000000000;//addi
//		ram[68] = 32'b00101000101001110000000000101011;//lw
//		ram[69] = 32'b00000100111010000000000000001101;//addi
//		ram[70] = 32'b00101001000001000000000000000000;//lw
//		ram[71] = 32'b00000100100111000000000000000000;//addi
//		ram[72] = 32'b00101000101001110000000000101011;//lw
//		ram[73] = 32'b00000100111010000000000000001110;//addi
//		ram[74] = 32'b00101001000001000000000000000000;//lw
//		ram[75] = 32'b00000100100111010000000000000000;//addi
//		ram[76] = 32'b00101000101001110000000000101011;//lw
//		ram[77] = 32'b00000100111010000000000000001111;//addi
//		ram[78] = 32'b00101001000001000000000000000000;//lw
//		ram[79] = 32'b00000100100111100000000000000000;//addi
//		ram[80] = 32'b00101000011111110000000000000001;//lw
//		ram[81] = 32'b00000011111000000000000000001100;//jr
//		ram[82] = 32'b00101100011111110000000000000001;//sw
//		ram[83] = 32'b00000100010000100000000000000001;//addi
//		ram[84] = 32'b00000100010000100000000000000001;//addi
//		ram[85] = 32'b00101000101001110000000000011011;//lw
//		ram[86] = 32'b00101000011010000000000000000010;//lw
//		ram[87] = 32'b00000000111010000100100000000001;//add
//		ram[88] = 32'b00101001001001110000000000000000;//lw
//		ram[89] = 32'b00101100101001110000000000101011;//sw
//		ram[90] = 32'b00000110000001000000000000000000;//addi
//		ram[91] = 32'b00101000101001110000000000101011;//lw
//		ram[92] = 32'b00101100111001000000000000000000;//sw
//		ram[93] = 32'b00000110001001000000000000000000;//addi
//		ram[94] = 32'b00101000101001110000000000101011;//lw
//		ram[95] = 32'b00000100111010000000000000000010;//addi
//		ram[96] = 32'b00101101000001000000000000000000;//sw
//		ram[97] = 32'b00000110010001000000000000000000;//addi
//		ram[98] = 32'b00101000101001110000000000101011;//lw
//		ram[99] = 32'b00000100111010000000000000000011;//addi
//		ram[100] = 32'b00101101000001000000000000000000;//sw
//		ram[101] = 32'b00000110011001000000000000000000;//addi
//		ram[102] = 32'b00101000101001110000000000101011;//lw
//		ram[103] = 32'b00000100111010000000000000000100;//addi
//		ram[104] = 32'b00101101000001000000000000000000;//sw
//		ram[105] = 32'b00000110100001000000000000000000;//addi
//		ram[106] = 32'b00101000101001110000000000101011;//lw
//		ram[107] = 32'b00000100111010000000000000000101;//addi
//		ram[108] = 32'b00101101000001000000000000000000;//sw
//		ram[109] = 32'b00000110101001000000000000000000;//addi
//		ram[110] = 32'b00101000101001110000000000101011;//lw
//		ram[111] = 32'b00000100111010000000000000000110;//addi
//		ram[112] = 32'b00101101000001000000000000000000;//sw
//		ram[113] = 32'b00000110110001000000000000000000;//addi
//		ram[114] = 32'b00101000101001110000000000101011;//lw
//		ram[115] = 32'b00000100111010000000000000000111;//addi
//		ram[116] = 32'b00101101000001000000000000000000;//sw
//		ram[117] = 32'b00000110111001000000000000000000;//addi
//		ram[118] = 32'b00101000101001110000000000101011;//lw
//		ram[119] = 32'b00000100111010000000000000001000;//addi
//		ram[120] = 32'b00101101000001000000000000000000;//sw
//		ram[121] = 32'b00000111000001000000000000000000;//addi
//		ram[122] = 32'b00101000101001110000000000101011;//lw
//		ram[123] = 32'b00000100111010000000000000001001;//addi
//		ram[124] = 32'b00101101000001000000000000000000;//sw
//		ram[125] = 32'b00000111001001000000000000000000;//addi
//		ram[126] = 32'b00101000101001110000000000101011;//lw
//		ram[127] = 32'b00000100111010000000000000001010;//addi
//		ram[128] = 32'b00101101000001000000000000000000;//sw
//		ram[129] = 32'b00000111010001000000000000000000;//addi
//		ram[130] = 32'b00101000101001110000000000101011;//lw
//		ram[131] = 32'b00000100111010000000000000001011;//addi
//		ram[132] = 32'b00101101000001000000000000000000;//sw
//		ram[133] = 32'b00000111011001000000000000000000;//addi
//		ram[134] = 32'b00101000101001110000000000101011;//lw
//		ram[135] = 32'b00000100111010000000000000001100;//addi
//		ram[136] = 32'b00101101000001000000000000000000;//sw
//		ram[137] = 32'b00000111100001000000000000000000;//addi
//		ram[138] = 32'b00101000101001110000000000101011;//lw
//		ram[139] = 32'b00000100111010000000000000001101;//addi
//		ram[140] = 32'b00101101000001000000000000000000;//sw
//		ram[141] = 32'b00000111101001000000000000000000;//addi
//		ram[142] = 32'b00101000101001110000000000101011;//lw
//		ram[143] = 32'b00000100111010000000000000001110;//addi
//		ram[144] = 32'b00101101000001000000000000000000;//sw
//		ram[145] = 32'b00000111110001000000000000000000;//addi
//		ram[146] = 32'b00101000101001110000000000101011;//lw
//		ram[147] = 32'b00000100111010000000000000001111;//addi
//		ram[148] = 32'b00101101000001000000000000000000;//sw
//		ram[149] = 32'b00101000011111110000000000000001;//lw
//		ram[150] = 32'b00000011111000000000000000001100;//jr
//		ram[151] = 32'b00000100000011110000000000000000;//addi
//		ram[152] = 32'b10010001111000000000000000000000;//show_pid
//		ram[153] = 32'b00101000101001110000000000010001;//lw
//		ram[154] = 32'b01100100111010000000000000000000;//seti
//		ram[155] = 32'b00011101000000000000000000010000;//beqz
//		ram[156] = 32'b00000100000011110000000000000000;//addi
//		ram[157] = 32'b00101100101011110000000000010000;//sw
//		ram[158] = 32'b00000100000011110000000000000001;//addi
//		ram[159] = 32'b00101100101011110000000000010001;//sw
//		ram[160] = 32'b00101000101001110000000000011111;//lw
//		ram[161] = 32'b00000100111010000000000000000000;//addi
//		ram[162] = 32'b00000100000011110000010000000000;//addi
//		ram[163] = 32'b00101101000011110000000000000000;//sw
//		ram[164] = 32'b00101000101001110000000000011111;//lw
//		ram[165] = 32'b00000100111010000000000000000001;//addi
//		ram[166] = 32'b00000100000011110000010100000000;//addi
//		ram[167] = 32'b00101101000011110000000000000000;//sw
//		ram[168] = 32'b00101000101001110000000000011111;//lw
//		ram[169] = 32'b00000100111010000000000000000010;//addi
//		ram[170] = 32'b00000100000011110000011000000000;//addi
//		ram[171] = 32'b00101101000011110000000000000000;//sw
//		ram[172] = 32'b00101000101001110000000000010000;//lw
//		ram[173] = 32'b01011000111010000000000000000000;//sgti
//		ram[174] = 32'b00011101000000000000000010000011;//beqz
//		ram[175] = 32'b00101000101001110000000000101100;//lw
//		ram[176] = 32'b01100100111010000000000000000001;//seti
//		ram[177] = 32'b00011101000000000000000000101100;//beqz
//		ram[178] = 32'b01101100100000000000000000000000;//get_pc
//		ram[179] = 32'b00101000101001110000000000010011;//lw
//		ram[180] = 32'b00101000101010000000000000010010;//lw
//		ram[181] = 32'b00000000111010000100100000000001;//add
//		ram[182] = 32'b00101101001001000000000000000000;//sw
//		ram[183] = 32'b00000111111001000000000000000000;//addi
//		ram[184] = 32'b00101100101001000000000000101110;//sw
//		ram[185] = 32'b00000110000001000000000000000000;//addi
//		ram[186] = 32'b00101000101001110000000000100011;//lw
//		ram[187] = 32'b00101000101010000000000000010010;//lw
//		ram[188] = 32'b00000000111010000100100000000001;//add
//		ram[189] = 32'b00101101001001000000000000000000;//sw
//		ram[190] = 32'b00101000101001110000000000100011;//lw
//		ram[191] = 32'b00101000101010000000000000010010;//lw
//		ram[192] = 32'b00000000111010000100100000000001;//add
//		ram[193] = 32'b00101001001001110000000000000000;//lw
//		ram[194] = 32'b01100100111010000000000000000000;//seti
//		ram[195] = 32'b00011101000000000000000000000100;//beqz
//		ram[196] = 32'b00101000101001110000000000010000;//lw
//		ram[197] = 32'b00000100111010001111111111111111;//addi
//		ram[198] = 32'b00101100101010000000000000010000;//sw
//		ram[199] = 32'b10001100110000000000000011011101;//jump_reg
//		ram[200] = 32'b00101000101001110000000000011011;//lw
//		ram[201] = 32'b00101000101010000000000000010010;//lw
//		ram[202] = 32'b00000000111010000100100000000001;//add
//		ram[203] = 32'b00101001001001110000000000000000;//lw
//		ram[204] = 32'b00000100111010000000000000000001;//addi
//		ram[205] = 32'b00101100101010000000000000101011;//sw
//		ram[206] = 32'b00101000101001110000000000101110;//lw
//		ram[207] = 32'b00101000101010000000000000101011;//lw
//		ram[208] = 32'b00101101000001110000000000000000;//sw
//		ram[209] = 32'b00101000101001110000000000010010;//lw
//		ram[210] = 32'b00101100010001110000000000000000;//sw
//		ram[211] = 32'b00000100010000100000000000000001;//addi
//		ram[212] = 32'b00101100010000110000000000000000;//sw
//		ram[213] = 32'b00000100010000110000000000000000;//addi
//		ram[214] = 32'b00000100010000100000000000000001;//addi
//		ram[215] = 32'b00101100011001110000000000000010;//sw
//		ram[216] = 32'b10001000110000000000000001010010;//jal_reg
//		ram[217] = 32'b00000100011000100000000000000000;//addi
//		ram[218] = 32'b00101000011000110000000000000000;//lw
//		ram[219] = 32'b00000100010000101111111111111111;//addi
//		ram[220] = 32'b00101000010001110000000000000000;//lw
//		ram[221] = 32'b10001100110000000000000011100110;//jump_reg
//		ram[222] = 32'b00101000101001110000000000100011;//lw
//		ram[223] = 32'b00101000101010000000000000010010;//lw
//		ram[224] = 32'b00000000111010000100100000000001;//add
//		ram[225] = 32'b00000100000011110000000000000000;//addi
//		ram[226] = 32'b00101101001011110000000000000000;//sw
//		ram[227] = 32'b00101000101001110000000000010000;//lw
//		ram[228] = 32'b00000100111010001111111111111111;//addi
//		ram[229] = 32'b00101100101010000000000000010000;//sw
//		ram[230] = 32'b00101000101001110000000000010000;//lw
//		ram[231] = 32'b01011000111010000000000000000000;//sgti
//		ram[232] = 32'b00011101000000000000000001000110;//beqz
//		ram[233] = 32'b00101000101001110000000000010010;//lw
//		ram[234] = 32'b00000100111010000000000000000001;//addi
//		ram[235] = 32'b00101100101010000000000000010010;//sw
//		ram[236] = 32'b00101000101001110000000000010010;//lw
//		ram[237] = 32'b01100100111010000000000000000011;//seti
//		ram[238] = 32'b00011101000000000000000000000010;//beqz
//		ram[239] = 32'b00000100000011110000000000000000;//addi
//		ram[240] = 32'b00101100101011110000000000010010;//sw
//		ram[241] = 32'b00101000101001110000000000100011;//lw
//		ram[242] = 32'b00101000101010000000000000010010;//lw
//		ram[243] = 32'b00000000111010000100100000000001;//add
//		ram[244] = 32'b00101001001001110000000000000000;//lw
//		ram[245] = 32'b01101000111010000000000000000001;//sdti
//		ram[246] = 32'b00011101000000000000000000001001;//beqz
//		ram[247] = 32'b00101000101001110000000000010010;//lw
//		ram[248] = 32'b00000100111010000000000000000001;//addi
//		ram[249] = 32'b00101100101010000000000000010010;//sw
//		ram[250] = 32'b00101000101001110000000000010010;//lw
//		ram[251] = 32'b01100100111010000000000000000011;//seti
//		ram[252] = 32'b00011101000000000000000000000010;//beqz
//		ram[253] = 32'b00000100000011110000000000000000;//addi
//		ram[254] = 32'b00101100101011110000000000010010;//sw
//		ram[255] = 32'b10001100110000000000000011110001;//jump_reg
//		ram[256] = 32'b00101000101001110000000000010010;//lw
//		ram[257] = 32'b00101100010001110000000000000000;//sw
//		ram[258] = 32'b00000100010000100000000000000001;//addi
//		ram[259] = 32'b00101100010000110000000000000000;//sw
//		ram[260] = 32'b00000100010000110000000000000000;//addi
//		ram[261] = 32'b00000100010000100000000000000001;//addi
//		ram[262] = 32'b00101100011001110000000000000010;//sw
//		ram[263] = 32'b10001000110000000000000000001101;//jal_reg
//		ram[264] = 32'b00000100011000100000000000000000;//addi
//		ram[265] = 32'b00101000011000110000000000000000;//lw
//		ram[266] = 32'b00000100010000101111111111111111;//addi
//		ram[267] = 32'b00101000010001110000000000000000;//lw
//		ram[268] = 32'b00101000101001110000000000011011;//lw
//		ram[269] = 32'b00101000101010000000000000010010;//lw
//		ram[270] = 32'b00000000111010000100100000000001;//add
//		ram[271] = 32'b00101001001001110000000000000000;//lw
//		ram[272] = 32'b00000100111010000000000000000001;//addi
//		ram[273] = 32'b00101100101010000000000000101011;//sw
//		ram[274] = 32'b00101000101001110000000000101011;//lw
//		ram[275] = 32'b00101000111001000000000000000000;//lw
//		ram[276] = 32'b00101100101001000000000000101010;//sw
//		ram[277] = 32'b00101000101001110000000000101010;//lw
//		ram[278] = 32'b00000100111111110000000000000000;//addi
//		ram[279] = 32'b00101000101001110000000000010000;//lw
//		ram[280] = 32'b01100100111010000000000000000001;//seti
//		ram[281] = 32'b00011101000000000000000000000010;//beqz
//		ram[282] = 32'b00000100000011110000000000000000;//addi
//		ram[283] = 32'b00101100101011110000000000101100;//sw
//		ram[284] = 32'b00101000101001110000000000010010;//lw
//		ram[285] = 32'b00000100111010000000000000000001;//addi
//		ram[286] = 32'b10010001000000000000000000000000;//show_pid
//		ram[287] = 32'b00101000101001110000000000101100;//lw
//		ram[288] = 32'b01100100111010000000000000000001;//seti
//		ram[289] = 32'b00011101000000000000000000000111;//beqz
//		ram[290] = 32'b00101000101001110000000000010011;//lw
//		ram[291] = 32'b00101000101010000000000000010010;//lw
//		ram[292] = 32'b00000000111010000100100000000001;//add
//		ram[293] = 32'b00101001001001110000000000000000;//lw
//		ram[294] = 32'b01110000000000000000000000000000;//enable_timer
//		ram[295] = 32'b00000000111000000000000000001100;//jr
//		ram[296] = 32'b10001100110000000000000100101110;//jump_reg
//		ram[297] = 32'b00101000101001110000000000010011;//lw
//		ram[298] = 32'b00101000101010000000000000010010;//lw
//		ram[299] = 32'b00000000111010000100100000000001;//add
//		ram[300] = 32'b00101001001001110000000000000000;//lw
//		ram[301] = 32'b00000000111000000000000000001100;//jr
//		ram[302] = 32'b10001100110000000000000100110001;//jump_reg
//		ram[303] = 32'b00000100000011110000001111100111;//addi
//		ram[304] = 32'b01010001111000000000000000000000;//output
//		ram[305] = 32'b10001100110000000000000111000010;//jump_reg
//		ram[306] = 32'b00000100000011110000000000000010;//addi
//		ram[307] = 32'b00101100101011110000000000010000;//sw
//		ram[308] = 32'b00000100000011110000000000000001;//addi
//		ram[309] = 32'b00101100101011110000000000101100;//sw
//		ram[310] = 32'b00000100000011110000000000000000;//addi
//		ram[311] = 32'b00101100101011110000000000101000;//sw
//		ram[312] = 32'b00101000101001110000000000101000;//lw
//		ram[313] = 32'b00101000101010000000000000010000;//lw
//		ram[314] = 32'b00000000111010000100100000001000;//slt
//		ram[315] = 32'b00011101001000000000000001011110;//beqz
//		ram[316] = 32'b00101000101001110000000000011111;//lw
//		ram[317] = 32'b00101000101010000000000000101000;//lw
//		ram[318] = 32'b00000000111010000100100000000001;//add
//		ram[319] = 32'b00101001001001110000000000000000;//lw
//		ram[320] = 32'b00101000101010000000000000010111;//lw
//		ram[321] = 32'b00101000101010010000000000101000;//lw
//		ram[322] = 32'b00000001000010010101000000000001;//add
//		ram[323] = 32'b00101101010001110000000000000000;//sw
//		ram[324] = 32'b00101000101001110000000000101000;//lw
//		ram[325] = 32'b00000100111010000000000000000001;//addi
//		ram[326] = 32'b00001001000001110000001000000000;//multi
//		ram[327] = 32'b00101000101010000000000000011011;//lw
//		ram[328] = 32'b00101000101010010000000000101000;//lw
//		ram[329] = 32'b00000001000010010101000000000001;//add
//		ram[330] = 32'b00101101010001110000000000000000;//sw
//		ram[331] = 32'b00101000101001110000000000011111;//lw
//		ram[332] = 32'b00101000101010000000000000101000;//lw
//		ram[333] = 32'b00000000111010000100100000000001;//add
//		ram[334] = 32'b00101001001001110000000000000000;//lw
//		ram[335] = 32'b00101000101010000000000000010011;//lw
//		ram[336] = 32'b00101000101010010000000000101000;//lw
//		ram[337] = 32'b00000001000010010101000000000001;//add
//		ram[338] = 32'b00101101010001110000000000000000;//sw
//		ram[339] = 32'b00101000101001110000000000100011;//lw
//		ram[340] = 32'b00101000101010000000000000101000;//lw
//		ram[341] = 32'b00000000111010000100100000000001;//add
//		ram[342] = 32'b00000100000011110000000000000001;//addi
//		ram[343] = 32'b00101101001011110000000000000000;//sw
//		ram[344] = 32'b00101000101001110000000000011011;//lw
//		ram[345] = 32'b00101000101010000000000000101000;//lw
//		ram[346] = 32'b00000000111010000100100000000001;//add
//		ram[347] = 32'b00101001001001110000000000000000;//lw
//		ram[348] = 32'b00000100111010000000000001000010;//addi
//		ram[349] = 32'b00101100101010000000000000101010;//sw
//		ram[350] = 32'b00101000101001110000000000011011;//lw
//		ram[351] = 32'b00101000101010000000000000101000;//lw
//		ram[352] = 32'b00000000111010000100100000000001;//add
//		ram[353] = 32'b00101001001001110000000000000000;//lw
//		ram[354] = 32'b00000100111010000000000000000010;//addi
//		ram[355] = 32'b00101100101010000000000000101011;//sw
//		ram[356] = 32'b00101000101001110000000000101010;//lw
//		ram[357] = 32'b00101000101010000000000000101011;//lw
//		ram[358] = 32'b00101101000001110000000000000000;//sw
//		ram[359] = 32'b00101000101001110000000000011011;//lw
//		ram[360] = 32'b00101000101010000000000000101000;//lw
//		ram[361] = 32'b00000000111010000100100000000001;//add
//		ram[362] = 32'b00101001001001110000000000000000;//lw
//		ram[363] = 32'b00000100111010000000000000000011;//addi
//		ram[364] = 32'b00101100101010000000000000101011;//sw
//		ram[365] = 32'b00101000101001110000000000101010;//lw
//		ram[366] = 32'b00101000101010000000000000101011;//lw
//		ram[367] = 32'b00101101000001110000000000000000;//sw
//		ram[368] = 32'b00101000101001110000000000011011;//lw
//		ram[369] = 32'b00101000101010000000000000101000;//lw
//		ram[370] = 32'b00000000111010000100100000000001;//add
//		ram[371] = 32'b00101001001001110000000000000000;//lw
//		ram[372] = 32'b00000100111010000000000000000101;//addi
//		ram[373] = 32'b00101100101010000000000000101011;//sw
//		ram[374] = 32'b00101000101001110000000000011011;//lw
//		ram[375] = 32'b00101000101010000000000000101000;//lw
//		ram[376] = 32'b00000000111010000100100000000001;//add
//		ram[377] = 32'b00101001001001110000000000000000;//lw
//		ram[378] = 32'b00101100101001110000000000101010;//sw
//		ram[379] = 32'b00101000101001110000000000101010;//lw
//		ram[380] = 32'b00101000101010000000000000101011;//lw
//		ram[381] = 32'b00101101000001110000000000000000;//sw
//		ram[382] = 32'b00101000101001110000000000011011;//lw
//		ram[383] = 32'b00101000101010000000000000101000;//lw
//		ram[384] = 32'b00000000111010000100100000000001;//add
//		ram[385] = 32'b00101001001001110000000000000000;//lw
//		ram[386] = 32'b00101100101001110000000000101011;//sw
//		ram[387] = 32'b00000100000011110000000000000001;//addi
//		ram[388] = 32'b00101100101011110000000000101010;//sw
//		ram[389] = 32'b00101000101001110000000000101010;//lw
//		ram[390] = 32'b00101000101010000000000000101011;//lw
//		ram[391] = 32'b00101101000001110000000000000000;//sw
//		ram[392] = 32'b00101000101001110000000000011011;//lw
//		ram[393] = 32'b00101000101010000000000000101000;//lw
//		ram[394] = 32'b00000000111010000100100000000001;//add
//		ram[395] = 32'b00101001001001110000000000000000;//lw
//		ram[396] = 32'b00000100111010000000000000000110;//addi
//		ram[397] = 32'b00101100101010000000000000101011;//sw
//		ram[398] = 32'b00101000101001110000000000010111;//lw
//		ram[399] = 32'b00101000101010000000000000101000;//lw
//		ram[400] = 32'b00000000111010000100100000000001;//add
//		ram[401] = 32'b00101001001001110000000000000000;//lw
//		ram[402] = 32'b00101100101001110000000000101010;//sw
//		ram[403] = 32'b00101000101001110000000000101010;//lw
//		ram[404] = 32'b00101000101010000000000000101011;//lw
//		ram[405] = 32'b00101101000001110000000000000000;//sw
//		ram[406] = 32'b00101000101001110000000000101000;//lw
//		ram[407] = 32'b00000100111010000000000000000001;//addi
//		ram[408] = 32'b00101100101010000000000000101000;//sw
//		ram[409] = 32'b10001100110000000000000100111000;//jump_reg
//		ram[410] = 32'b00000100000011110000000000000000;//addi
//		ram[411] = 32'b00101100101011110000000000010010;//sw
//		ram[412] = 32'b00101100010000110000000000000000;//sw
//		ram[413] = 32'b00000100010000110000000000000000;//addi
//		ram[414] = 32'b00000100010000100000000000000001;//addi
//		ram[415] = 32'b00000100000011110000000000000000;//addi
//		ram[416] = 32'b00101100011011110000000000000010;//sw
//		ram[417] = 32'b10001000110000000000000000001101;//jal_reg
//		ram[418] = 32'b00000100011000100000000000000000;//addi
//		ram[419] = 32'b00101000011000110000000000000000;//lw
//		ram[420] = 32'b00101000101001110000000000011011;//lw
//		ram[421] = 32'b00000100111010000000000000000000;//addi
//		ram[422] = 32'b00101001000001110000000000000000;//lw
//		ram[423] = 32'b00000100111010000000000000000001;//addi
//		ram[424] = 32'b00101100101010000000000000101011;//sw
//		ram[425] = 32'b00101000101001110000000000101011;//lw
//		ram[426] = 32'b00101000111001000000000000000000;//lw
//		ram[427] = 32'b00101100101001000000000000101010;//sw
//		ram[428] = 32'b00101000101001110000000000101010;//lw
//		ram[429] = 32'b00000100111111110000000000000000;//addi
//		ram[430] = 32'b00101000101001110000000000010000;//lw
//		ram[431] = 32'b01100100111010000000000000000001;//seti
//		ram[432] = 32'b00011101000000000000000000000010;//beqz
//		ram[433] = 32'b00000100000011110000000000000000;//addi
//		ram[434] = 32'b00101100101011110000000000101100;//sw
//		ram[435] = 32'b00000100000011110000000000000001;//addi
//		ram[436] = 32'b10010001111000000000000000000000;//show_pid
//		ram[437] = 32'b00101000101001110000000000101100;//lw
//		ram[438] = 32'b01100100111010000000000000000001;//seti
//		ram[439] = 32'b00011101000000000000000000000110;//beqz
//		ram[440] = 32'b00101000101001110000000000010011;//lw
//		ram[441] = 32'b00000100111010000000000000000000;//addi
//		ram[442] = 32'b00101001000001110000000000000000;//lw
//		ram[443] = 32'b01110000000000000000000000000000;//enable_timer
//		ram[444] = 32'b00000000111000000000000000001100;//jr
//		ram[445] = 32'b10001100110000000000000111000010;//jump_reg
//		ram[446] = 32'b00101000101001110000000000010011;//lw
//		ram[447] = 32'b00000100111010000000000000000000;//addi
//		ram[448] = 32'b00101001000001110000000000000000;//lw
//		ram[449] = 32'b00000000111000000000000000001100;//jr



//		ram[1024] = 32'b01000100000000000000000000000000;//nop
//		ram[1025] = 32'b01000100000000000000000000000000;//nop
//		ram[1026] = 32'b10001110101000000000000000000011;//jump_reg
//		ram[1027] = 32'b00000110001100010000000000000001;//addi
//		ram[1028] = 32'b00000100000101100000000000000111;//addi
//		ram[1029] = 32'b00000110110101101111111111111001;//addi
//		ram[1030] = 32'b00101110010101100000000000000000;//sw
//		ram[1031] = 32'b00000100000100000000000000000000;//addi
//		ram[1032] = 32'b01110100000000000000000000000000;//disable_timer
//		ram[1033] = 32'b00111100000000000000000010010111;//jump

		ram[1024] = 32'b01000100000000000000000000000000;//nop
		ram[1025] = 32'b01000100000000000000000000000000;//nop
		ram[1026] = 32'b10001110101000000000000000000011;//jump_reg
		ram[1027] = 32'b00000110001100010000000000000001;//addi
		ram[1028] = 32'b00000100000101100000000000000111;//addi
		ram[1029] = 32'b00000110110101101111111111111001;//addi
		ram[1030] = 32'b00101110010101100000000000000000;//sw
		ram[1031] = 32'b00101010010101100000000000000000;//lw
		ram[1032] = 32'b01010010110000000000000000000000;//output
		ram[1033] = 32'b00000100000100000000000000000000;//addi
		ram[1034] = 32'b01110100000000000000000000000000;//disable_timer
		ram[1035] = 32'b00111100000000000000000010010111;//jump

		
//		ram[1280] = 32'b01000100000000000000000000000000;//nop
//		ram[1281] = 32'b01000100000000000000000000000000;//nop
//		ram[1282] = 32'b10001110101000000000000000000011;//jump_reg
//		ram[1283] = 32'b00000110001100010000000000000001;//addi
//		ram[1284] = 32'b00000100000101100000000000000111;//addi
//		ram[1285] = 32'b00001010110101100000000000000111;//multi
//		ram[1286] = 32'b00101110010101100000000000000000;//sw
//		ram[1287] = 32'b00000100000100000000000000000000;//addi
//		ram[1288] = 32'b01110100000000000000000000000000;//disable_timer
//		ram[1289] = 32'b00111100000000000000000010010111;//jump

		ram[1280] = 32'b01000100000000000000000000000000;//nop
		ram[1281] = 32'b01000100000000000000000000000000;//nop
		ram[1282] = 32'b10001110101000000000000000000011;//jump_reg
		ram[1283] = 32'b00000110001100010000000000000001;//addi
		ram[1284] = 32'b00000100000101100000000000000111;//addi
		ram[1285] = 32'b00001010110101100000000000000111;//multi
		ram[1286] = 32'b00101110010101100000000000000000;//sw
		ram[1287] = 32'b00101010010101100000000000000000;//lw
		ram[1288] = 32'b01010010110000000000000000000000;//output
		ram[1289] = 32'b00000100000100000000000000000000;//addi
		ram[1290] = 32'b01110100000000000000000000000000;//disable_timer
		ram[1291] = 32'b00111100000000000000000010010111;//jump
		
//		ram[1536] = 32'b01000100000000000000000000000000;//nop
//		ram[1537] = 32'b01000100000000000000000000000000;//nop
//		ram[1538] = 32'b10001110101000000000000000000011;//jump_reg
//		ram[1539] = 32'b00000110001100010000000000000001;//addi
//		ram[1540] = 32'b00000100000101100000000000000111;//addi
//		ram[1541] = 32'b00001110110101100000000000000111;//divi
//		ram[1542] = 32'b00101110010101100000000000000000;//sw
//		ram[1543] = 32'b00101010010101100000000000000000;//lw
//		ram[1544] = 32'b01010010110000000000000000000000;//output
//		ram[1545] = 32'b00000100000100000000000000000000;//addi
//		ram[1546] = 32'b01110100000000000000000000000000;//disable_timer
//		ram[1547] = 32'b00111100000000000000000010010111;//jump

		ram[1536] = 32'b01000100000000000000000000000000;//nop
		ram[1537] = 32'b01000100000000000000000000000000;//nop
		ram[1538] = 32'b10001110101000000000000000000011;//jump_reg
		ram[1539] = 32'b00000110001100010000000000000001;//addi
		ram[1540] = 32'b00000100000101100000000000000111;//addi
		ram[1541] = 32'b00001110110101100000000000000111;//divi
		ram[1542] = 32'b00101110010101100000000000000000;//sw
		ram[1543] = 32'b00000100000100000000000000000000;//addi
		ram[1544] = 32'b01110100000000000000000000000000;//disable_timer
		ram[1545] = 32'b00111100000000000000000010010111;//jump





	end 
	
	
	always @ (posedge write_clock)
	begin
		// Write
		if (we)
			ram[write_addr] <= data;
	end
	
	always @ (posedge read_clock)
	begin
		// Read 
		q <= ram[read_addr];
	end
	
endmodule
